module top_module(output out, input in);
  assign out=~in;
endmodule
